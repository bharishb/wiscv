`define FIXED_LATENCY
`define SYNTHESIS
`define FPGA_MODE